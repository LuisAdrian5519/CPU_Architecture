-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: User
-- 
-- Create Date:    06/06/2024 01:22:12
-- Project Name:   Procesador
-- Module Name:    Procesador.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Procesador is
    port(
        X: in std_logic_vector(8 downto 0);
        SalALU: out std_logic_vector(8 downto 0);
--        Oper: in std_logic_vector(4 downto 0); --debseria ser se;al
        Cout: out std_logic;
        CLK: in std_logic;
--        MUX1, MUX2: in std_logic_vector(1 downto 0);se;al
        Instr: out std_logic_vector(8 downto 0);
--        address: in std_logic_vector(8 downto 0);--no port
        data_out: out std_logic_vector(15 downto 0);
         Dout: out std_logic_vector(8 downto 0)
    );
end Procesador;

architecture arq1 of Procesador is
    signal R1, R2, R3: std_logic_vector(8 downto 0) := "000000000";
    signal OUT1, OUT2: std_logic_vector(8 downto 0);
    signal ALU_result_with_carry: std_logic_vector(9 downto 0);--?
    signal R: std_logic_vector(8 downto 0);
    signal CLRPC, INCPC, LDMAR, LDMBR, LDIR, OEPC, LDPC, OEMBR, OEALU, RD, WR, LDR1, LDR2, LDR3: std_logic := '0';
    signal PCOut, BusDir, BusDatos, MBROut, BUSD0, BUSD1: std_logic_vector(8 downto 0) := "000000000";
    signal InstrReg: std_logic_vector(8 downto 0) := (others => '0');
    signal Scontrol: std_logic_vector(15 downto 0);
    signal WR_signal, RD_signal, LDR1_signal, LDR2_signal, LDR3_signal: std_logic;
    type RAM_type is array (0 to 2423) of std_logic_vector(15 downto 0);
	signal Oper: std_logic_vector(4 downto 0);
	signal MUX1, MUX2: std_logic_vector(1 downto 0);
    signal RAM_content: RAM_type := (
--000 NOP
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 	
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000",x"0000", x"0000", 
--010 SUM
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",--SUM R1, #
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",--SUM R1, R1
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",--SUM R1, R2
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",--SUM R1, R3
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",--SUM R2, #
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",--SUM R2, R1
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",--SUM R2, R2
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",--SUM R2, R3
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",--SUM R3, #
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",--SUM R3, R1     
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",--SUM R3, R2
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000", --SUM R3, R3
--020 SUB
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

--030 MUL
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
		x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

--040 DIV
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
		
--050 COMPLEMENTO
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0029", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0025", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0023", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",

--060 AND
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

--070 OR
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

-- 080 XOR
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

--090 SHR
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",

--0A0 SHL
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",

--0B0 INC
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",

-- 0C0 DEC
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",

-- 0D0 MOV
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

-- 0E0 CMP
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0003", x"0000", x"0000", x"0000", x"0000",

-- 180 MOV Memoria - Registro
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0820", x"1040", x"0029",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0029", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0820", x"1040", x"0025",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0025", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0820", x"1040", x"0023",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0023", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0801", x"1040", x"0023", x"0000", x"0000",

-- 190 MOV Registro - Memoria
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0820", x"0041", x"2020",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0820", x"0041", x"2020",
	x"0B00", x"1040", x"0030", x"0B00", x"1040", x"0820", x"0041", x"2020",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",
	x"0B00", x"1040", x"0030", x"0041", x"0820", x"0041", x"2020", x"0000",

-- 100 RD
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"1009", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"1005", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"1003", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",

-- 110 WR
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0400", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000",
	x"0B00", x"1040", x"0030", x"0000", x"0000", x"0000", x"0000", x"0000"


      
    );
    signal paso: std_logic_vector(2 downto 0) := "000";
    signal a: std_logic_vector(11 downto 0);
    type Mem_RAM is array (0 to 3) of std_logic_vector(8 downto 0);
    signal contenido : Mem_RAM := ( 
        "011010001", -- MOV R1, X
        "011001001", -- MOV R2, R1 (calcular 2x)
        "011011001", -- MOV R3, #1
        "000011001"  -- SUM R2, R1 (sumar 2x y 1)
    );
begin
    SalALU <= R;

    Reg1: process(LDR1, CLK)
    variable tmp1: std_logic_vector(8 downto 0) := "000000000";
    begin
        if rising_edge(CLK) and LDR1 = '1' then
            tmp1 := R;
        end if;
        R1 <= tmp1;
    end process;

    Reg2: process(LDR2, CLK)
    variable tmp2: std_logic_vector(8 downto 0) := "000000000";
    begin
        if rising_edge(CLK) and LDR2 = '1' then
            tmp2 := R;
        end if;
        R2 <= tmp2;
    end process;

    Reg3: process(LDR3, CLK)
    variable tmp3: std_logic_vector(8 downto 0) := "000000000";
    begin
        if rising_edge(CLK) and LDR3 = '1' then
            tmp3 := R;
        end if;
        R3 <= tmp3;
    end process;

    process(MUX1, MUX2, BUSD0, R1, R2, R3)
    begin
        case MUX1 is
            when "00" => OUT1 <= BUSD0;
            when "01" => OUT1 <= R1;
            when "10" => OUT1 <= R2;
            when "11" => OUT1 <= R3;
            when others => OUT1 <= "000000000";
        end case;

        case MUX2 is
            when "00" => OUT2 <= BUSD0;
            when "01" => OUT2 <= R1;
            when "10" => OUT2 <= R2;
            when "11" => OUT2 <= R3;
            when others => OUT2 <= "000000000";
        end case;
    end process;

    process (Oper, OUT1, OUT2)
    variable At, Bt, Rt: std_logic_vector(9 downto 0);
    begin
        At := '0' & OUT1;
        Bt := '0' & OUT2;
        case Oper is
            when "00000" =>
                Rt := At;
                Cout <= '0';
            when "00001" =>
                Rt := std_logic_vector(unsigned(At) + unsigned(Bt));
                Cout <= Rt(9);
            when others =>
                Rt := "ZZZZZZZZZZ";
        end case;
        ALU_result_with_carry <= Rt;
        R <= Rt(8 downto 0);
    end process;

    PC: process(CLRPC, INCPC, CLK, OEPC, LDPC, BUSD0)
    variable tmp: std_logic_vector(8 downto 0) := "000000000";
    begin
        if rising_edge(CLK) then
            if CLRPC = '1' then
                tmp := "000000000";
            elsif INCPC = '1' then
                tmp := std_logic_vector(unsigned(tmp) + 1);
            end if;
        end if;
        if OEPC = '1' then 
            BUSD0 <= tmp;
        else 
            BUSD0 <= "ZZZZZZZZZ";
        end if;
    end process;

    MAR: process(LDMAR, CLK, PCout, BUSD0)
    variable tmp: std_logic_vector(8 downto 0) := "000000000";
    begin
        if rising_edge(CLK) and LDMAR = '1' then
            tmp := BUSD0;
        end if;
        BusDir <= tmp;
    end process;

    MBR: process(LDMBR, CLK, BUSD1, OEMBR)
    variable tmp: std_logic_vector(8 downto 0) := "000000000";
    begin
        if rising_edge(CLK) and LDMBR = '1' then
            tmp := BUSD1;
        end if;
		if OEMBR ='0' then
		BUSD0 <= "ZZZZZZZZZ";
		else
		BUSD0 <= tmp;
		end if;
--debe tener 3er estado
    end process;

    IR: process(LDIR, CLK, BUSD0)
    variable tmp: std_logic_vector(8 downto 0) := (others => '0');
    begin
---weird
        if rising_edge(CLK) and LDIR = '1' then
            tmp := BUSD0;
        end if;
        InstrReg <= tmp;
        Instr <= InstrReg;
    end process;

    WR <= Scontrol(13);
    RD <= Scontrol(12);
    LDMAR <= Scontrol(11);
    CLRPC <= Scontrol(10);
    INCPC <= Scontrol(9);
    OEPC <= Scontrol(8);
    LDPC <= Scontrol(7);
    LDMBR <= Scontrol(6);
    OEMBR <= Scontrol(5);
    LDIR <= Scontrol(4);
    LDR1_signal <= Scontrol(3);
    LDR2_signal <= Scontrol(2);
    LDR3_signal <= Scontrol(1);
    OEALU <= Scontrol(0);
	Oper <= InstrReg(8 downto 4);
	MUX1 <= InstrReg(3 downto 2);
	MUX2 <= InstrReg(1 downto 0);

    process(clk)
    begin
--        a <= address & paso;
			a <= InstrReg & paso;
        if rising_edge(clk) then
            paso <= std_logic_vector(unsigned(paso) + 1);
--            data_out <= RAM_content(to_integer(unsigned(a)));
        end if;
				data_out <= RAM_content(to_integer(unsigned(a)));
    end process;

    process(BUSDir, BUSD0, rd, wr, clk)
    variable palabra: integer range 0 to 7;
    begin
        palabra := to_integer(unsigned(BUSDir));
        if rising_edge(clk) then
            if rd = '1' then
                BUSD1 <= contenido(palabra);
            elsif wr = '1' then
                contenido(palabra) <= BUSD0;
                BUSD1 <= (others => 'Z');
            else
                BUSD1 <= (others => 'Z');
            end if;
        end if;
    end process;
end arq1;


