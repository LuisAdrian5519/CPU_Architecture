-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: User
-- 
-- Create Date:    15/03/2024 02:02:53
-- Project Name:   Compemento1
-- Module Name:    Compemento1.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity Compemento1 is
--   port( );
end Compemento1;

architecture arq1 of Compemento1 is
begin

end arq1;
